*Design
vin in 0 pulse (0 2.101 100p 50p 50p 200p 500p)
r1 in out 1.01k
c1 out 0 101f

*Stimulation
.tran 20ps 1500ps

*Plotting
.control
run
set color0=white
plot v(in),v(out)
set hcopydevtype=postscript
hardcopy rc1.ps v(out) v(in) 
.endc
.end
