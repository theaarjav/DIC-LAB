*TTL Inverter vtc

.model transistor npn Q(BF=20.2)
Vcc vcc 0 5v
Vin ip 0 5v

Q1 b b1 ip transistor
Q2 op b 0 transistor
Rc vcc op 1.01k
Rb vcc b1 10k

.DC vin 0 5 0.01
.control
run
set color0=white
set color1=black
plot v(vout)
set hcopydevtype=postscript
hardcopy rc1.ps v(vout)
.endc
.end


.DC vin 0 5 0.01
.control
run
set color0=white
plot v(op)
set hcopydevtype=postscript
hardcopy rc1.ps v(op)
.endc
.end
