*TTL Inverter

Q1 b b1 ip transistor
Q2 op b 0 transistor
Rc vcc op 1.01k
Rb vcc b1 10.1k
Vcc vcc 0 5v
Vin ip 0 pulse (0 5 120p 10p 10p 150p 400p)

.tran 1ps 400ps

.control
run
set color0=white
plot v(op) v(ip)
set hcopydevtype=postscript
hardcopy rc1.ps v(op)
.endc
.end
.model transistor npn Q(BF=20.2)