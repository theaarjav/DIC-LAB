magic
tech scmos
timestamp 1681066144
<< nwell >>
rect -18 1 20 18
<< polysilicon >>
rect -8 8 -6 11
rect 8 8 10 11
rect -8 -2 -6 3
rect 8 -2 10 3
rect -8 -12 -6 -6
rect 8 -12 10 -6
rect -8 -20 -6 -16
rect 8 -20 10 -16
<< ndiffusion >>
rect -12 -16 -8 -12
rect -6 -16 8 -12
rect 10 -16 14 -12
<< pdiffusion >>
rect -12 3 -8 8
rect -6 3 8 8
rect 10 3 14 8
<< metal1 >>
rect -16 8 -12 12
rect 14 -2 18 3
rect -4 -6 -2 -2
rect 4 -6 6 -2
rect 14 -6 22 -2
rect 14 -12 18 -6
rect -16 -20 -12 -16
<< ntransistor >>
rect -8 -16 -6 -12
rect 8 -16 10 -12
<< ptransistor >>
rect -8 3 -6 8
rect 8 3 10 8
<< polycontact >>
rect -8 -6 -4 -2
rect 6 -6 10 -2
<< ndcontact >>
rect -16 -16 -12 -12
rect 14 -16 18 -12
<< pdcontact >>
rect -16 3 -12 8
rect 14 3 18 8
<< psubstratepcontact >>
rect -16 -24 -12 -20
<< nsubstratencontact >>
rect -16 12 -12 16
<< labels >>
rlabel nsubstratencontact -16 16 -12 16 4 vdd_101
rlabel psubstratepcontact -16 -24 -12 -24 2 gnd
rlabel metal1 -2 -6 -2 -2 1 va_101
rlabel metal1 4 -6 4 -2 1 vb_101
rlabel metal1 22 -6 22 -2 7 vout_101
<< end >>
