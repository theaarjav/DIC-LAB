magic
tech scmos
timestamp 1681040728
<< nwell >>
rect -22 2 18 20
<< polysilicon >>
rect -12 10 -10 13
rect 6 10 8 13
rect -12 -6 -10 3
rect 6 -6 8 3
rect -12 -13 -10 -10
rect 6 -13 8 -10
rect -12 -21 -10 -17
rect 6 -21 8 -17
<< ndiffusion >>
rect -16 -17 -12 -13
rect -10 -17 6 -13
rect 8 -17 12 -13
<< pdiffusion >>
rect -20 9 -12 10
rect -16 5 -12 9
rect -20 3 -12 5
rect -10 9 6 10
rect -10 5 -4 9
rect 0 5 6 9
rect -10 3 6 5
rect 8 9 16 10
rect 8 5 12 9
rect 8 3 16 5
<< metal1 >>
rect -20 14 -4 18
rect 0 14 16 18
rect -20 9 -16 14
rect 12 9 16 14
rect -4 1 0 5
rect -24 -3 0 1
rect -20 -13 -16 -3
rect -8 -10 -6 -6
rect 10 -10 12 -6
rect 12 -21 16 -17
<< ntransistor >>
rect -12 -17 -10 -13
rect 6 -17 8 -13
<< ptransistor >>
rect -12 3 -10 10
rect 6 3 8 10
<< polycontact >>
rect -12 -10 -8 -6
rect 6 -10 10 -6
<< ndcontact >>
rect -20 -17 -16 -13
rect 12 -17 16 -13
<< pdcontact >>
rect -20 5 -16 9
rect -4 5 0 9
rect 12 5 16 9
<< psubstratepcontact >>
rect 12 -25 16 -21
<< nsubstratencontact >>
rect -4 14 0 18
<< labels >>
rlabel psubstratepcontact 12 -25 16 -25 8 gnd_96
rlabel metal1 -24 -3 -24 1 3 vout_96
rlabel nsubstratencontact -4 18 0 18 5 vdd_96
rlabel metal1 12 -10 12 -6 1 vb_96
rlabel metal1 -6 -10 -6 -6 1 va_96
<< end >>
