*CMOS Circuit
.include cmos_90nm.txt

vdd d1 0 1.2v
*vgs g1 0 pulse(0 1.2v 20ns 0ns 0ns 180ns 500ns)
vgs g1 0 1.2v

.subckt fanout d1 g1 0 out 
M1 d1 g1 out d1 PMOS w=5u l=0.09u
M2 out g1 0 0  NMOS w=1u l=0.09u
.ends fanout

x d1 g1 0 out fanout
c1 out 0 10pf
x1 d1 out 0 out1 fanout
x2 d1 out 0 out2 fanout
x3 d1 out 0 out3 fanout
x4 d1 out 0 out4 fanout
x5 d1 out 0 out5 fanout
x6 d1 out 0 out6 fanout
x7 d1 out 0 out7 fanout
x8 d1 out 0 out8 fanout
x9 d1 out 0 out9 fanout
x10 d1 out 0 out10 fanout
x11 d1 out 0 out11 fanout
x12 d1 out 0 out12 fanout
x13 d1 out 0 out13 fanout
x14 d1 out 0 out14 fanout
x15 d1 out 0 out15 fanout
x16 d1 out 0 out16 fanout
x17 d1 out 0 out17 fanout
x18 d1 out 0 out18 fanout
x19 d1 out 0 out19 fanout
x20 d1 out 0 out20 fanout


.control
*tran 1ns 1000ns
dc vgs 0 1.2v 0.01

plot v(out), v(g1)
.endc
.end
