*Design
Va va 0 pulse (0 5 120p 10p 10p 150p 400p)
 Vb vb 0 pulse (0 5 120p 10p 10p 440p 900p)
 Vcc vcc 0 5v

Q1a b2 b1 va transistor 
Q1b b2 b1 vb transistor 
Q2 c2 b2 e2 transistor 
Q3 vcc c2 vout transistor 
Q4 vout e2 0 transistor 
Rb1 vcc b1 10.1k
Rc1 vcc c2 1.01k
 Rc2 c2 0 10.1k

.tran 1ps 1000ps

.control 
Run
Set color0=white
plot v(vout) 
plot v(vb) v(va)
set hcopydevtype=postscript
 hardcopy rc1.ps v(vout)
.endc
.end
.model transistor npn Q(BF=20.2)
